package my_testbench_pkg;
  import uvm_pkg::*;

//============================================================
// 1.  Declare distinct IMP types
//============================================================
`uvm_analysis_imp_decl(_exp)
`uvm_analysis_imp_decl(_act)

//============================================================
// 2.  Simple transaction
//============================================================
class my_txn extends uvm_sequence_item;
  rand int data;
  `uvm_object_utils(my_txn)
  function new(string name="my_txn"); super.new(name); endfunction
  function string convert2string(); return $sformatf("data=%0d", data); endfunction
endclass

//============================================================
// 3.  Producers: two simple monitors
//============================================================
class exp_monitor extends uvm_component;
  `uvm_component_utils(exp_monitor)
  uvm_analysis_port #(my_txn) ap;
  function new(string name, uvm_component parent); super.new(name,parent); endfunction
  function void build_phase(uvm_phase phase); ap = new("ap", this); endfunction
  task run_phase(uvm_phase phase);
    my_txn t;
    repeat (5) begin
      t = my_txn::type_id::create("t");
      t.randomize() with { data inside {[0:9]}; }; // expected stream
      ap.write(t);
      #5ns;
    end
  endtask
endclass

class act_monitor extends uvm_component;
  `uvm_component_utils(act_monitor)
  uvm_analysis_port #(my_txn) ap;
  function new(string name, uvm_component parent); super.new(name,parent); endfunction
  function void build_phase(uvm_phase phase); ap = new("ap", this); endfunction
  task run_phase(uvm_phase phase);
    my_txn t;
    repeat (5) begin
      t = my_txn::type_id::create("t");
      t.randomize() with { data inside {[0:9]}; }; // actual stream
      ap.write(t);
      #7ns;
    end
  endtask
endclass

//============================================================
// 4.  Scoreboard with TWO imps
//============================================================
class my_scoreboard extends uvm_component;
  `uvm_component_utils(my_scoreboard)

  // create two imps with unique suffixes
  uvm_analysis_imp_exp #(my_txn, my_scoreboard) exp_imp;
  uvm_analysis_imp_act #(my_txn, my_scoreboard) act_imp;

  // Queues to hold incoming txns
  my_txn exp_q[$], act_q[$];

  function new(string name, uvm_component parent); super.new(name,parent); endfunction

  function void build_phase(uvm_phase phase);
    exp_imp = new("exp_imp", this);
    act_imp = new("act_imp", this);
  endfunction

  // These are generated by the IMP typedefs:
  //   function void write_exp(my_txn t);
  //   function void write_act(my_txn t);
  function void write_exp(my_txn t);
    `uvm_info("SCOREBOARD", $sformatf("EXP got %s", t.convert2string()), UVM_LOW)
    exp_q.push_back(t);
    compare_if_ready();
  endfunction

  function void write_act(my_txn t);
    `uvm_info("SCOREBOARD", $sformatf("ACT got %s", t.convert2string()), UVM_LOW)
    act_q.push_back(t);
    compare_if_ready();
  endfunction

  function void compare_if_ready();
    if (exp_q.size() && act_q.size()) begin
      my_txn e = exp_q.pop_front();
      my_txn a = act_q.pop_front();
      if (e.data == a.data)
        `uvm_info("SCOREBOARD", $sformatf("MATCH  exp=%0d act=%0d", e.data, a.data), UVM_MEDIUM)
      else
        `uvm_error("SCOREBOARD", $sformatf("MISMATCH exp=%0d act=%0d", e.data, a.data))
    end
  endfunction
endclass
  
 class my_env extends uvm_env;
  `uvm_component_utils(my_env)
  exp_monitor     m_exp_mon;
  act_monitor     m_act_mon;
  my_scoreboard   m_scb;

  function new(string name, uvm_component parent); super.new(name,parent); endfunction

  function void build_phase(uvm_phase phase);
    m_exp_mon = exp_monitor   ::type_id::create("m_exp_mon", this);
    m_act_mon = act_monitor   ::type_id::create("m_act_mon", this);
    m_scb     = my_scoreboard ::type_id::create("m_scb",     this);
  endfunction

  function void connect_phase(uvm_phase phase);
    m_exp_mon.ap.connect(m_scb.exp_imp);
    m_act_mon.ap.connect(m_scb.act_imp);
  endfunction
endclass
  
class my_test extends uvm_test;
  `uvm_component_utils(my_test)
  my_env m_env;
  function new(string name, uvm_component parent); super.new(name,parent); endfunction
  function void build_phase(uvm_phase phase);
    m_env = my_env::type_id::create("m_env", this);
  endfunction
endclass
  
endpackage